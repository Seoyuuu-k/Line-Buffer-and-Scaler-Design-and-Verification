`include "top.v"
`include "single_port_ram.v"
`include "video_timing.sv" 